// miniProject.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module miniProject (
		input  wire        clk_clk,            //         clk.clk
		output wire [10:0] lcd_wire_export,    //    lcd_wire.export
		output wire [9:0]  led_wire_export,    //    led_wire.export
		output wire [3:0]  motor_wire_export,  //  motor_wire.export
		input  wire        reset_reset,        //       reset.reset
		output wire        sdram_clk_clk,      //   sdram_clk.clk
		output wire [12:0] sdram_wire_addr,    //  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,      //            .ba
		output wire        sdram_wire_cas_n,   //            .cas_n
		output wire        sdram_wire_cke,     //            .cke
		output wire        sdram_wire_cs_n,    //            .cs_n
		inout  wire [15:0] sdram_wire_dq,      //            .dq
		output wire [1:0]  sdram_wire_dqm,     //            .dqm
		output wire        sdram_wire_ras_n,   //            .ras_n
		output wire        sdram_wire_we_n,    //            .we_n
		input  wire [9:0]  switch_wire_export  // switch_wire.export
	);

	wire         sys_sdram_pll_0_sys_clk_clk;                                 // sys_sdram_pll_0:sys_clk_clk -> [CPU:clk, DMEM:clk, LCD:clk, LED:clk, MEMORY:clk, MOTOR:clk, SWITCH:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, rst_controller:clk, rst_controller_001:clk, sysid_qsys_0:clock, timer_0:clk, timer_1:clk]
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                                 // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                     // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                  // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                        // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_readdatavalid;                               // mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	wire         cpu_data_master_write;                                       // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                   // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                              // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                 // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                        // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;              // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;           // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;           // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;               // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                  // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;            // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                 // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;             // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                      // mm_interconnect_0:MEMORY_s1_chipselect -> MEMORY:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                        // MEMORY:readdata -> mm_interconnect_0:MEMORY_s1_readdata
	wire  [15:0] mm_interconnect_0_memory_s1_address;                         // mm_interconnect_0:MEMORY_s1_address -> MEMORY:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                      // mm_interconnect_0:MEMORY_s1_byteenable -> MEMORY:byteenable
	wire         mm_interconnect_0_memory_s1_write;                           // mm_interconnect_0:MEMORY_s1_write -> MEMORY:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                       // mm_interconnect_0:MEMORY_s1_writedata -> MEMORY:writedata
	wire         mm_interconnect_0_memory_s1_clken;                           // mm_interconnect_0:MEMORY_s1_clken -> MEMORY:clken
	wire         mm_interconnect_0_dmem_s1_chipselect;                        // mm_interconnect_0:DMEM_s1_chipselect -> DMEM:az_cs
	wire  [15:0] mm_interconnect_0_dmem_s1_readdata;                          // DMEM:za_data -> mm_interconnect_0:DMEM_s1_readdata
	wire         mm_interconnect_0_dmem_s1_waitrequest;                       // DMEM:za_waitrequest -> mm_interconnect_0:DMEM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_dmem_s1_address;                           // mm_interconnect_0:DMEM_s1_address -> DMEM:az_addr
	wire         mm_interconnect_0_dmem_s1_read;                              // mm_interconnect_0:DMEM_s1_read -> DMEM:az_rd_n
	wire   [1:0] mm_interconnect_0_dmem_s1_byteenable;                        // mm_interconnect_0:DMEM_s1_byteenable -> DMEM:az_be_n
	wire         mm_interconnect_0_dmem_s1_readdatavalid;                     // DMEM:za_valid -> mm_interconnect_0:DMEM_s1_readdatavalid
	wire         mm_interconnect_0_dmem_s1_write;                             // mm_interconnect_0:DMEM_s1_write -> DMEM:az_wr_n
	wire  [15:0] mm_interconnect_0_dmem_s1_writedata;                         // mm_interconnect_0:DMEM_s1_writedata -> DMEM:az_data
	wire         mm_interconnect_0_lcd_s1_chipselect;                         // mm_interconnect_0:LCD_s1_chipselect -> LCD:chipselect
	wire  [31:0] mm_interconnect_0_lcd_s1_readdata;                           // LCD:readdata -> mm_interconnect_0:LCD_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_s1_address;                            // mm_interconnect_0:LCD_s1_address -> LCD:address
	wire         mm_interconnect_0_lcd_s1_write;                              // mm_interconnect_0:LCD_s1_write -> LCD:write_n
	wire  [31:0] mm_interconnect_0_lcd_s1_writedata;                          // mm_interconnect_0:LCD_s1_writedata -> LCD:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                         // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                           // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                            // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_write;                              // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                          // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                        // SWITCH:readdata -> mm_interconnect_0:SWITCH_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                         // mm_interconnect_0:SWITCH_s1_address -> SWITCH:address
	wire         mm_interconnect_0_motor_s1_chipselect;                       // mm_interconnect_0:MOTOR_s1_chipselect -> MOTOR:chipselect
	wire  [31:0] mm_interconnect_0_motor_s1_readdata;                         // MOTOR:readdata -> mm_interconnect_0:MOTOR_s1_readdata
	wire   [1:0] mm_interconnect_0_motor_s1_address;                          // mm_interconnect_0:MOTOR_s1_address -> MOTOR:address
	wire         mm_interconnect_0_motor_s1_write;                            // mm_interconnect_0:MOTOR_s1_write -> MOTOR:write_n
	wire  [31:0] mm_interconnect_0_motor_s1_writedata;                        // mm_interconnect_0:MOTOR_s1_writedata -> MOTOR:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver0_irq;                                    // timer_1:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                                 // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [CPU:reset_n, DMEM:reset_n, MEMORY:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, timer_0:reset_n, timer_1:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [CPU:reset_req, MEMORY:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                               // CPU:debug_reset_request -> rst_controller:reset_in0
	wire         sys_sdram_pll_0_reset_source_reset;                          // sys_sdram_pll_0:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [LCD:reset_n, LED:reset_n, MOTOR:reset_n, SWITCH:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, sysid_qsys_0:reset_n]

	miniProject_CPU cpu (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                       //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	miniProject_DMEM dmem (
		.clk            (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),         // reset.reset_n
		.az_addr        (mm_interconnect_0_dmem_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_dmem_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_dmem_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_dmem_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_dmem_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_dmem_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_dmem_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_dmem_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_dmem_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                         //  wire.export
		.zs_ba          (sdram_wire_ba),                           //      .export
		.zs_cas_n       (sdram_wire_cas_n),                        //      .export
		.zs_cke         (sdram_wire_cke),                          //      .export
		.zs_cs_n        (sdram_wire_cs_n),                         //      .export
		.zs_dq          (sdram_wire_dq),                           //      .export
		.zs_dqm         (sdram_wire_dqm),                          //      .export
		.zs_ras_n       (sdram_wire_ras_n),                        //      .export
		.zs_we_n        (sdram_wire_we_n)                          //      .export
	);

	miniProject_LCD lcd (
		.clk        (sys_sdram_pll_0_sys_clk_clk),         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_lcd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_s1_readdata),   //                    .readdata
		.out_port   (lcd_wire_export)                      // external_connection.export
	);

	miniProject_LED led (
		.clk        (sys_sdram_pll_0_sys_clk_clk),         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_wire_export)                      // external_connection.export
	);

	miniProject_MEMORY memory (
		.clk        (sys_sdram_pll_0_sys_clk_clk),            //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	miniProject_MOTOR motor (
		.clk        (sys_sdram_pll_0_sys_clk_clk),           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_motor_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_motor_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_motor_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_motor_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_motor_s1_readdata),   //                    .readdata
		.out_port   (motor_wire_export)                      // external_connection.export
	);

	miniProject_SWITCH switch (
		.clk      (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_wire_export)                    // external_connection.export
	);

	miniProject_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	miniProject_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                        //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_0_reset_source_reset)  // reset_source.reset
	);

	miniProject_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_sdram_pll_0_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	miniProject_timer_0 timer_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	miniProject_timer_0 timer_1 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	miniProject_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_0_sys_clk_clk                   (sys_sdram_pll_0_sys_clk_clk),                                 //                 sys_sdram_pll_0_sys_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                              //         CPU_reset_reset_bridge_in_reset.reset
		.jtag_uart_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // jtag_uart_0_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                       (cpu_data_master_address),                                     //                         CPU_data_master.address
		.CPU_data_master_waitrequest                   (cpu_data_master_waitrequest),                                 //                                        .waitrequest
		.CPU_data_master_byteenable                    (cpu_data_master_byteenable),                                  //                                        .byteenable
		.CPU_data_master_read                          (cpu_data_master_read),                                        //                                        .read
		.CPU_data_master_readdata                      (cpu_data_master_readdata),                                    //                                        .readdata
		.CPU_data_master_readdatavalid                 (cpu_data_master_readdatavalid),                               //                                        .readdatavalid
		.CPU_data_master_write                         (cpu_data_master_write),                                       //                                        .write
		.CPU_data_master_writedata                     (cpu_data_master_writedata),                                   //                                        .writedata
		.CPU_data_master_debugaccess                   (cpu_data_master_debugaccess),                                 //                                        .debugaccess
		.CPU_instruction_master_address                (cpu_instruction_master_address),                              //                  CPU_instruction_master.address
		.CPU_instruction_master_waitrequest            (cpu_instruction_master_waitrequest),                          //                                        .waitrequest
		.CPU_instruction_master_read                   (cpu_instruction_master_read),                                 //                                        .read
		.CPU_instruction_master_readdata               (cpu_instruction_master_readdata),                             //                                        .readdata
		.CPU_instruction_master_readdatavalid          (cpu_instruction_master_readdatavalid),                        //                                        .readdatavalid
		.CPU_debug_mem_slave_address                   (mm_interconnect_0_cpu_debug_mem_slave_address),               //                     CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write                     (mm_interconnect_0_cpu_debug_mem_slave_write),                 //                                        .write
		.CPU_debug_mem_slave_read                      (mm_interconnect_0_cpu_debug_mem_slave_read),                  //                                        .read
		.CPU_debug_mem_slave_readdata                  (mm_interconnect_0_cpu_debug_mem_slave_readdata),              //                                        .readdata
		.CPU_debug_mem_slave_writedata                 (mm_interconnect_0_cpu_debug_mem_slave_writedata),             //                                        .writedata
		.CPU_debug_mem_slave_byteenable                (mm_interconnect_0_cpu_debug_mem_slave_byteenable),            //                                        .byteenable
		.CPU_debug_mem_slave_waitrequest               (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),           //                                        .waitrequest
		.CPU_debug_mem_slave_debugaccess               (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),           //                                        .debugaccess
		.DMEM_s1_address                               (mm_interconnect_0_dmem_s1_address),                           //                                 DMEM_s1.address
		.DMEM_s1_write                                 (mm_interconnect_0_dmem_s1_write),                             //                                        .write
		.DMEM_s1_read                                  (mm_interconnect_0_dmem_s1_read),                              //                                        .read
		.DMEM_s1_readdata                              (mm_interconnect_0_dmem_s1_readdata),                          //                                        .readdata
		.DMEM_s1_writedata                             (mm_interconnect_0_dmem_s1_writedata),                         //                                        .writedata
		.DMEM_s1_byteenable                            (mm_interconnect_0_dmem_s1_byteenable),                        //                                        .byteenable
		.DMEM_s1_readdatavalid                         (mm_interconnect_0_dmem_s1_readdatavalid),                     //                                        .readdatavalid
		.DMEM_s1_waitrequest                           (mm_interconnect_0_dmem_s1_waitrequest),                       //                                        .waitrequest
		.DMEM_s1_chipselect                            (mm_interconnect_0_dmem_s1_chipselect),                        //                                        .chipselect
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.LCD_s1_address                                (mm_interconnect_0_lcd_s1_address),                            //                                  LCD_s1.address
		.LCD_s1_write                                  (mm_interconnect_0_lcd_s1_write),                              //                                        .write
		.LCD_s1_readdata                               (mm_interconnect_0_lcd_s1_readdata),                           //                                        .readdata
		.LCD_s1_writedata                              (mm_interconnect_0_lcd_s1_writedata),                          //                                        .writedata
		.LCD_s1_chipselect                             (mm_interconnect_0_lcd_s1_chipselect),                         //                                        .chipselect
		.LED_s1_address                                (mm_interconnect_0_led_s1_address),                            //                                  LED_s1.address
		.LED_s1_write                                  (mm_interconnect_0_led_s1_write),                              //                                        .write
		.LED_s1_readdata                               (mm_interconnect_0_led_s1_readdata),                           //                                        .readdata
		.LED_s1_writedata                              (mm_interconnect_0_led_s1_writedata),                          //                                        .writedata
		.LED_s1_chipselect                             (mm_interconnect_0_led_s1_chipselect),                         //                                        .chipselect
		.MEMORY_s1_address                             (mm_interconnect_0_memory_s1_address),                         //                               MEMORY_s1.address
		.MEMORY_s1_write                               (mm_interconnect_0_memory_s1_write),                           //                                        .write
		.MEMORY_s1_readdata                            (mm_interconnect_0_memory_s1_readdata),                        //                                        .readdata
		.MEMORY_s1_writedata                           (mm_interconnect_0_memory_s1_writedata),                       //                                        .writedata
		.MEMORY_s1_byteenable                          (mm_interconnect_0_memory_s1_byteenable),                      //                                        .byteenable
		.MEMORY_s1_chipselect                          (mm_interconnect_0_memory_s1_chipselect),                      //                                        .chipselect
		.MEMORY_s1_clken                               (mm_interconnect_0_memory_s1_clken),                           //                                        .clken
		.MOTOR_s1_address                              (mm_interconnect_0_motor_s1_address),                          //                                MOTOR_s1.address
		.MOTOR_s1_write                                (mm_interconnect_0_motor_s1_write),                            //                                        .write
		.MOTOR_s1_readdata                             (mm_interconnect_0_motor_s1_readdata),                         //                                        .readdata
		.MOTOR_s1_writedata                            (mm_interconnect_0_motor_s1_writedata),                        //                                        .writedata
		.MOTOR_s1_chipselect                           (mm_interconnect_0_motor_s1_chipselect),                       //                                        .chipselect
		.SWITCH_s1_address                             (mm_interconnect_0_switch_s1_address),                         //                               SWITCH_s1.address
		.SWITCH_s1_readdata                            (mm_interconnect_0_switch_s1_readdata),                        //                                        .readdata
		.sysid_qsys_0_control_slave_address            (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //              sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata           (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                        .readdata
		.timer_0_s1_address                            (mm_interconnect_0_timer_0_s1_address),                        //                              timer_0_s1.address
		.timer_0_s1_write                              (mm_interconnect_0_timer_0_s1_write),                          //                                        .write
		.timer_0_s1_readdata                           (mm_interconnect_0_timer_0_s1_readdata),                       //                                        .readdata
		.timer_0_s1_writedata                          (mm_interconnect_0_timer_0_s1_writedata),                      //                                        .writedata
		.timer_0_s1_chipselect                         (mm_interconnect_0_timer_0_s1_chipselect),                     //                                        .chipselect
		.timer_1_s1_address                            (mm_interconnect_0_timer_1_s1_address),                        //                              timer_1_s1.address
		.timer_1_s1_write                              (mm_interconnect_0_timer_1_s1_write),                          //                                        .write
		.timer_1_s1_readdata                           (mm_interconnect_0_timer_1_s1_readdata),                       //                                        .readdata
		.timer_1_s1_writedata                          (mm_interconnect_0_timer_1_s1_writedata),                      //                                        .writedata
		.timer_1_s1_chipselect                         (mm_interconnect_0_timer_1_s1_chipselect)                      //                                        .chipselect
	);

	miniProject_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (sys_sdram_pll_0_reset_source_reset), // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
